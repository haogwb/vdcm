module xfm_rec #(parameter BPC=8)
(
input clk,
input rstn,

input [5:0] bpv2x2[0:3],
input [5:0] bpv2x1_p0[0:3],
input [5:0] bpv2x1_p1[0:3]
);


endmodule
