`timescale 1ns/1ps

module tb;

bit clk;

bit rstn;

initial begin

  forever #10ns clk = ~clk; 

end



initial begin

 rstn = 1'b0; 

 #20ns;

 rstn = 1'b1; 

 #32us;

 //$stop;
 $finish;

end



bit [127:0] codec_data;
bit [127:0] codec_data_ssm1;
bit [127:0] codec_data_ssm2;
bit [127:0] codec_data_ssm3;

bit codec_data_rd_en;
bit codec_data_rd_en_ssm1;
bit codec_data_rd_en_ssm2;
bit codec_data_rd_en_ssm3;
bit start_dec;
bit start_dec_ff;
bit start_dec_ff1;
initial begin
  #1us;
  @(posedge clk) start_dec <= 1;
//  @(posedge clk) start_dec_ff = 1;
//  @(posedge clk) start_dec_ff1 = 1;
end

always@(posedge clk)begin
  start_dec_ff <= start_dec;
  start_dec_ff1 <= start_dec_ff;
end
wire [10:0] blk_x;
wire [10:0] blk_y;
reg [9:0] c;
reg [9:0] r;
always@(posedge clk or negedge rstn)begin
  if(~rstn)
    c <= 'd0;
  else if(start_dec_ff1)
    if(c==1080/8-1)
       c <= 0;
    else
       c <= c+'d1;
end

always@(posedge clk or negedge rstn)begin
  if(~rstn)
    r <= 'd0;
  else if(start_dec_ff1)
    if(c==1080/8-1)
       r <= r+'d1;
end

assign blk_x = c*8;
assign blk_y = r*2;
wire isFls = r==0;
wire isNxtBlkFls = isFls & c<1080/8-1; 

wire [7:0] mpp_qres_ssm0 [0:16-1];
reg  [7:0] mpp_qres_ssm0_ff [0:16-1];
wire [7:0] mpp_qres_ssm1 [0:16-1];
wire [7:0] mpp_qres_ssm2 [0:16-1];
wire [7:0] mpp_qres_ssm3 [0:16-1];

wire modeNxt_XFM;
wire modeNxt_BP;
wire modeNxt_MPPF;
wire [3:0] use2x2;
wire [3:0] modeNxt_Mpp_stepsize;

wire [8:0]xfm_coeff_0 ; 
wire [8:0]xfm_coeff_1 ; 
wire [8:0]xfm_coeff_2 ; 
wire [8:0]xfm_coeff_3 ; 
wire [8:0]xfm_coeff_4 ; 
wire [8:0]xfm_coeff_5 ; 
wire [8:0]xfm_coeff_6 ; 
wire [8:0]xfm_coeff_7 ; 
wire [8:0]xfm_coeff_8 ; 
wire [8:0]xfm_coeff_9 ; 
wire [8:0]xfm_coeff_10; 
wire [8:0]xfm_coeff_11; 
wire [8:0]xfm_coeff_12; 
wire [8:0]xfm_coeff_13; 
wire [8:0]xfm_coeff_14; 
wire [8:0]xfm_coeff_15; 
bitparse #(.ssm_idx(0)) u_bitparse(

  .clk     (clk),

  .rstn     (rstn),
  .start_dec (start_dec),
  .codec_data_rd_en (codec_data_rd_en),

  .codec_data       (codec_data),
  .isNxtBlockFls    (isNxtBlkFls), 

  .modeNxt_XFM      (modeNxt_XFM),
  .modeNxt_BP       (modeNxt_BP),
  .modeNxt_MPPF       (modeNxt_MPPF),
  .use2x2           (use2x2),
  .modeNxt_Mpp_stepsize(modeNxt_Mpp_stepsize),
  .pnxtBlkQuant(mpp_qres_ssm0)

);
bitparse_ssm123 #(.ssm_idx(1)) u_bitparse_ssm1(

  .clk     (clk),

  .rstn     (rstn),
  .start_dec (start_dec_ff),
  .codec_data_rd_en (codec_data_rd_en_ssm1),

  .codec_data       (codec_data_ssm1),
  .isFls            (isFls),
  .modeNxt_XFM      (modeNxt_XFM),
  .modeNxt_BP       (modeNxt_BP),
  .modeNxt_MPPF       (modeNxt_MPPF),
  .use2x2           (use2x2[1]),
  .modeNxt_Mpp_stepsize(modeNxt_Mpp_stepsize),

  .pnxtBlkQuant(mpp_qres_ssm1),

  .xfm_coeff_0   (xfm_coeff_0 ) ,
  .xfm_coeff_1   (xfm_coeff_1 ) ,
  .xfm_coeff_2   (xfm_coeff_2 ) ,
  .xfm_coeff_3   (xfm_coeff_3 ) ,
  .xfm_coeff_4   (xfm_coeff_4 ) ,
  .xfm_coeff_5   (xfm_coeff_5 ) ,
  .xfm_coeff_6   (xfm_coeff_6 ) ,
  .xfm_coeff_7   (xfm_coeff_7 ) ,
  .xfm_coeff_8   (xfm_coeff_8 ) ,
  .xfm_coeff_9   (xfm_coeff_9 ) ,
  .xfm_coeff_10  (xfm_coeff_10) ,
  .xfm_coeff_11  (xfm_coeff_11) ,
  .xfm_coeff_12  (xfm_coeff_12) ,
  .xfm_coeff_13  (xfm_coeff_13) ,
  .xfm_coeff_14  (xfm_coeff_14) ,
  .xfm_coeff_15  (xfm_coeff_15) 
);
bitparse_ssm123 #(.ssm_idx(2)) u_bitparse_ssm2(

  .clk     (clk),

  .rstn     (rstn),
  .start_dec (start_dec_ff),
  .codec_data_rd_en (codec_data_rd_en_ssm2),

  .codec_data       (codec_data_ssm2),

  .isFls            (isFls),
  .modeNxt_XFM      (modeNxt_XFM),
  .modeNxt_BP       (modeNxt_BP),
  .modeNxt_MPPF       (modeNxt_MPPF),
  .use2x2           (use2x2[2]),
  .modeNxt_Mpp_stepsize(modeNxt_Mpp_stepsize),

  .pnxtBlkQuant(mpp_qres_ssm2)
);

bitparse_ssm123 #(.ssm_idx(3)) u_bitparse_ssm3(

  .clk     (clk),

  .rstn     (rstn),
  .start_dec (start_dec_ff),
  .codec_data_rd_en (codec_data_rd_en_ssm3),

  .codec_data       (codec_data_ssm3),

  .isFls            (isFls),
  .modeNxt_XFM      (modeNxt_XFM),
  .modeNxt_BP       (modeNxt_BP),
  .modeNxt_MPPF       (modeNxt_MPPF),
  .use2x2           (use2x2[3]),
  .modeNxt_Mpp_stepsize(modeNxt_Mpp_stepsize),

  .pnxtBlkQuant(mpp_qres_ssm3)
);

always@(posedge clk)
  mpp_qres_ssm0_ff <= mpp_qres_ssm0;
decMpp  u_decMpp (
    .clk     (clk),
    .rstn     (rstn),
    .blk_vld         ( start_dec_ff),
    .mpp_qres_ssm0   ( mpp_qres_ssm0_ff ),
    .mpp_qres_ssm1   ( mpp_qres_ssm1 ),
    .mpp_qres_ssm2   ( mpp_qres_ssm2 ),
    .mpp_qres_ssm3   ( mpp_qres_ssm3 )
);


xfm_rec  u_xfm_rec (
    .clk                     ( clk                 ),
    .rstn                    ( rstn                ),
    .coeff_0             ( xfm_coeff_0   [8:0] ),
    .coeff_1             ( xfm_coeff_1   [8:0] ),
    .coeff_2             ( xfm_coeff_2   [8:0] ),
    .coeff_3             ( xfm_coeff_3   [8:0] ),
    .coeff_4             ( xfm_coeff_4   [8:0] ),
    .coeff_5             ( xfm_coeff_5   [8:0] ),
    .coeff_6             ( xfm_coeff_6   [8:0] ),
    .coeff_7             ( xfm_coeff_7   [8:0] ),
    .coeff_8             ( xfm_coeff_8   [8:0] ),
    .coeff_9             ( xfm_coeff_9   [8:0] ),
    .coeff_10            ( xfm_coeff_10  [8:0] ),
    .coeff_11            ( xfm_coeff_11  [8:0] ),
    .coeff_12            ( xfm_coeff_12  [8:0] ),
    .coeff_13            ( xfm_coeff_13  [8:0] ),
    .coeff_14            ( xfm_coeff_14  [8:0] ),
    .coeff_15            ( xfm_coeff_15  [8:0] )
);


  

reg [127:0] codec_bits[0:4050-1];

initial begin

$readmemh("./bits.bits",codec_bits);

end



bit [10:0] codec_rd_addr;
bit [2:0] rd_en_num;
assign rd_en_num =  codec_data_rd_en + codec_data_rd_en_ssm1 + codec_data_rd_en_ssm2 + codec_data_rd_en_ssm3;
always@(posedge clk or negedge rstn)
  if(~rstn)
    codec_rd_addr <= 0;
  else if(rd_en_num==4)
    codec_rd_addr <= codec_rd_addr + 4;
  else if(rd_en_num==3)
    codec_rd_addr <= codec_rd_addr + 3;
  else if(rd_en_num==2)
    codec_rd_addr <= codec_rd_addr + 2;
  else if(rd_en_num==1)
    codec_rd_addr <= codec_rd_addr + 1;

always@(*)
begin
  if(codec_data_rd_en)
  codec_data = codec_bits[codec_rd_addr];

  if(codec_data_rd_en & codec_data_rd_en_ssm1)
    codec_data_ssm1 = codec_bits[codec_rd_addr+1];
  else if(codec_data_rd_en_ssm1)
    codec_data_ssm1 = codec_bits[codec_rd_addr];

  if(codec_data_rd_en & codec_data_rd_en_ssm1& codec_data_rd_en_ssm2)
    codec_data_ssm2 = codec_bits[codec_rd_addr+2];
  else if((codec_data_rd_en ^ codec_data_rd_en_ssm1)& codec_data_rd_en_ssm2)
    codec_data_ssm2 = codec_bits[codec_rd_addr+1];
  else if(codec_data_rd_en_ssm2)
    codec_data_ssm2 = codec_bits[codec_rd_addr+0];

  if(codec_data_rd_en & codec_data_rd_en_ssm1& codec_data_rd_en_ssm2& codec_data_rd_en_ssm3)
    codec_data_ssm3 = codec_bits[codec_rd_addr+3];
  else if((codec_data_rd_en+codec_data_rd_en_ssm1+ codec_data_rd_en_ssm2)==2 & codec_data_rd_en_ssm3)
    codec_data_ssm3 = codec_bits[codec_rd_addr+2];
  else if((codec_data_rd_en+codec_data_rd_en_ssm1+ codec_data_rd_en_ssm2)==1 & codec_data_rd_en_ssm3)
    codec_data_ssm3 = codec_bits[codec_rd_addr+1];
  else 
    codec_data_ssm3 = codec_bits[codec_rd_addr+0];


//  if(codec_data_rd_en)

//    codec_rd_addr = codec_rd_addr + 1;

end



initial begin

    $fsdbDumpfile("test.fsdb");

    $fsdbDumpvars(0,tb);

    $fsdbDumpMDA(0, tb);

end



endmodule;
