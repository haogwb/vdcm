module decVecEcSymbolSM #(parameter ssm_idx = 0)
(
input [127:0] suffix,
input [1:0] bitsReq,
output reg[7:0] symbol,
output reg[1:0] mask,
output [7:0] size,

output [8:0] src_0,
output [8:0] src_1,
output [8:0] src_2,
output [8:0] src_3
);


wire [2:0] vecGrk = 5;
wire [7:0] maxPrefix = ((1<<(bitsReq*4))-1) >>vecGrk;
wire [7:0] uiBits = suffix[127-:8];
reg [3:0] prefix_tmp;
always@(*)
begin
  prefix_tmp = 0;
  casez (uiBits)
    8'b0???_????: prefix_tmp = 0;
    8'b10??_????: prefix_tmp = 1;
    8'b110?_????: prefix_tmp = 2;
    8'b1110_????: prefix_tmp = 3;
    8'b1111_0???: prefix_tmp = 4;
    8'b1111_10??: prefix_tmp = 5;
    8'b1111_110?: prefix_tmp = 6;
    8'b1111_1110: prefix_tmp = 7;
    8'b1111_1111: prefix_tmp = 8;
    default:prefix_tmp = 0;
  endcase
end

wire [3:0] prefix = prefix_tmp > maxPrefix  ? maxPrefix : prefix_tmp;
wire [3:0] prefix_size = prefix+1;

wire [127:0] suffix_rm_prefix = suffix<<prefix_size;
wire [7:0] gf_suffix = suffix_rm_prefix[127-:5];//vecGrk];
wire [7:0] vecCodeNum = (prefix<<vecGrk) | gf_suffix;

wire [3:0] vec_sm_bitsReq_1_luma_inv [0:15];
wire [4-1:0] vec_sm_bitsReq_1_chroma_inv[0:15];
wire [8-1:0]vec_sm_bitsReq_2_luma_inv[0:255];
wire [8-1:0]vec_sm_bitsReq_2_chroma_inv[0:255]; 

always@(*)
begin
  case(bitsReq)
    2'd1: symbol = ssm_idx==1 ? vec_sm_bitsReq_1_luma_inv[vecCodeNum] : vec_sm_bitsReq_1_chroma_inv[vecCodeNum];
    2'd2: symbol = ssm_idx==1 ? vec_sm_bitsReq_2_luma_inv[vecCodeNum] : vec_sm_bitsReq_2_chroma_inv[vecCodeNum];
  endcase
end
always@(*)
begin
  case(bitsReq)
    2'd1: mask=1;
    2'd2: mask=3;
  endcase
end


wire [7:0] maxValue = (1<<bitsReq) -1;
assign src_0 = (symbol >> (bitsReq*3)) & mask;
assign src_1 = (symbol >> (bitsReq*2)) & mask;
assign src_2 = (symbol >> (bitsReq*1)) & mask;
assign src_3 = (symbol >> (bitsReq*0)) & mask;

assign size = prefix_size + vecGrk;


assign vec_sm_bitsReq_1_luma_inv[00] = 4'd2;
assign vec_sm_bitsReq_1_luma_inv[01] = 4'd1;
assign vec_sm_bitsReq_1_luma_inv[02] = 4'd8;
assign vec_sm_bitsReq_1_luma_inv[03] = 4'd4;
assign vec_sm_bitsReq_1_luma_inv[04] = 4'd10;
assign vec_sm_bitsReq_1_luma_inv[05] = 4'd5;
assign vec_sm_bitsReq_1_luma_inv[06] = 4'd3;
assign vec_sm_bitsReq_1_luma_inv[07] = 4'd9;
assign vec_sm_bitsReq_1_luma_inv[08] = 4'd6;
assign vec_sm_bitsReq_1_luma_inv[09] = 4'd12;
assign vec_sm_bitsReq_1_luma_inv[10] = 4'd7;
assign vec_sm_bitsReq_1_luma_inv[11] = 4'd11;
assign vec_sm_bitsReq_1_luma_inv[12] = 4'd14;
assign vec_sm_bitsReq_1_luma_inv[13] = 4'd13;
assign vec_sm_bitsReq_1_luma_inv[14] = 4'd15;
assign vec_sm_bitsReq_1_luma_inv[15] = 4'd0;

assign vec_sm_bitsReq_1_chroma_inv[0] = 2;
assign vec_sm_bitsReq_1_chroma_inv[1] = 1;
assign vec_sm_bitsReq_1_chroma_inv[2] = 4;
assign vec_sm_bitsReq_1_chroma_inv[3] = 8;
assign vec_sm_bitsReq_1_chroma_inv[4] = 3;
assign vec_sm_bitsReq_1_chroma_inv[5] = 12;
assign vec_sm_bitsReq_1_chroma_inv[6] = 10;
assign vec_sm_bitsReq_1_chroma_inv[7] = 5;
assign vec_sm_bitsReq_1_chroma_inv[8] = 6;
assign vec_sm_bitsReq_1_chroma_inv[9] = 9;
assign vec_sm_bitsReq_1_chroma_inv[10] = 11;
assign vec_sm_bitsReq_1_chroma_inv[11] = 7;
assign vec_sm_bitsReq_1_chroma_inv[12] = 13;
assign vec_sm_bitsReq_1_chroma_inv[13] = 14;
assign vec_sm_bitsReq_1_chroma_inv[14] = 15;
assign vec_sm_bitsReq_1_chroma_inv[15] = 0;


assign vec_sm_bitsReq_2_luma_inv[0] =8;
assign vec_sm_bitsReq_2_luma_inv[1] =2;
assign vec_sm_bitsReq_2_luma_inv[2] =128;
assign vec_sm_bitsReq_2_luma_inv[3] =32;
assign vec_sm_bitsReq_2_luma_inv[4] =6;
assign vec_sm_bitsReq_2_luma_inv[5] =9;
assign vec_sm_bitsReq_2_luma_inv[6] =18;
assign vec_sm_bitsReq_2_luma_inv[7] =72;
assign vec_sm_bitsReq_2_luma_inv[8] =132;
assign vec_sm_bitsReq_2_luma_inv[9] =33;
assign vec_sm_bitsReq_2_luma_inv[10] =66;
assign vec_sm_bitsReq_2_luma_inv[11] =24;
assign vec_sm_bitsReq_2_luma_inv[12] =129;
assign vec_sm_bitsReq_2_luma_inv[13] =36;
assign vec_sm_bitsReq_2_luma_inv[14] =144;
assign vec_sm_bitsReq_2_luma_inv[15] =96;
assign vec_sm_bitsReq_2_luma_inv[16] =22;
assign vec_sm_bitsReq_2_luma_inv[17] =73;
assign vec_sm_bitsReq_2_luma_inv[18] =12;
assign vec_sm_bitsReq_2_luma_inv[19] =3;
assign vec_sm_bitsReq_2_luma_inv[20] =25;
assign vec_sm_bitsReq_2_luma_inv[21] =70;
assign vec_sm_bitsReq_2_luma_inv[22] =88;
assign vec_sm_bitsReq_2_luma_inv[23] =82;
assign vec_sm_bitsReq_2_luma_inv[24] =37;
assign vec_sm_bitsReq_2_luma_inv[25] =133;
assign vec_sm_bitsReq_2_luma_inv[26] =148;
assign vec_sm_bitsReq_2_luma_inv[27] =97;
assign vec_sm_bitsReq_2_luma_inv[28] =192;
assign vec_sm_bitsReq_2_luma_inv[29] =48;
assign vec_sm_bitsReq_2_luma_inv[30] =145;
assign vec_sm_bitsReq_2_luma_inv[31] =100;
assign vec_sm_bitsReq_2_luma_inv[32] =86;
assign vec_sm_bitsReq_2_luma_inv[33] =89;
assign vec_sm_bitsReq_2_luma_inv[34] =10;
assign vec_sm_bitsReq_2_luma_inv[35] =34;
assign vec_sm_bitsReq_2_luma_inv[36] =136;
assign vec_sm_bitsReq_2_luma_inv[37] =149;
assign vec_sm_bitsReq_2_luma_inv[38] =101;
assign vec_sm_bitsReq_2_luma_inv[39] =13;
assign vec_sm_bitsReq_2_luma_inv[40] =7;
assign vec_sm_bitsReq_2_luma_inv[41] =76;
assign vec_sm_bitsReq_2_luma_inv[42] =19;
assign vec_sm_bitsReq_2_luma_inv[43] =160;
assign vec_sm_bitsReq_2_luma_inv[44] =40;
assign vec_sm_bitsReq_2_luma_inv[45] =49;
assign vec_sm_bitsReq_2_luma_inv[46] =28;
assign vec_sm_bitsReq_2_luma_inv[47] =67;
assign vec_sm_bitsReq_2_luma_inv[48] =130;
assign vec_sm_bitsReq_2_luma_inv[49] =196;
assign vec_sm_bitsReq_2_luma_inv[50] =112;
assign vec_sm_bitsReq_2_luma_inv[51] =208;
assign vec_sm_bitsReq_2_luma_inv[52] =52;
assign vec_sm_bitsReq_2_luma_inv[53] =193;
assign vec_sm_bitsReq_2_luma_inv[54] =74;
assign vec_sm_bitsReq_2_luma_inv[55] =38;
assign vec_sm_bitsReq_2_luma_inv[56] =26;
assign vec_sm_bitsReq_2_luma_inv[57] =137;
assign vec_sm_bitsReq_2_luma_inv[58] =98;
assign vec_sm_bitsReq_2_luma_inv[59] =152;
assign vec_sm_bitsReq_2_luma_inv[60] =77;
assign vec_sm_bitsReq_2_luma_inv[61] =41;
assign vec_sm_bitsReq_2_luma_inv[62] =23;
assign vec_sm_bitsReq_2_luma_inv[63] =83;
assign vec_sm_bitsReq_2_luma_inv[64] =71;
assign vec_sm_bitsReq_2_luma_inv[65] =29;
assign vec_sm_bitsReq_2_luma_inv[66] =92;
assign vec_sm_bitsReq_2_luma_inv[67] =90;
assign vec_sm_bitsReq_2_luma_inv[68] =134;
assign vec_sm_bitsReq_2_luma_inv[69] =164;
assign vec_sm_bitsReq_2_luma_inv[70] =153;
assign vec_sm_bitsReq_2_luma_inv[71] =146;
assign vec_sm_bitsReq_2_luma_inv[72] =104;
assign vec_sm_bitsReq_2_luma_inv[73] =161;
assign vec_sm_bitsReq_2_luma_inv[74] =113;
assign vec_sm_bitsReq_2_luma_inv[75] =102;
assign vec_sm_bitsReq_2_luma_inv[76] =53;
assign vec_sm_bitsReq_2_luma_inv[77] =197;
assign vec_sm_bitsReq_2_luma_inv[78] =212;
assign vec_sm_bitsReq_2_luma_inv[79] =209;
assign vec_sm_bitsReq_2_luma_inv[80] =116;
assign vec_sm_bitsReq_2_luma_inv[81] =165;
assign vec_sm_bitsReq_2_luma_inv[82] =14;
assign vec_sm_bitsReq_2_luma_inv[83] =150;
assign vec_sm_bitsReq_2_luma_inv[84] =11;
assign vec_sm_bitsReq_2_luma_inv[85] =35;
assign vec_sm_bitsReq_2_luma_inv[86] =93;
assign vec_sm_bitsReq_2_luma_inv[87] =105;
assign vec_sm_bitsReq_2_luma_inv[88] =50;
assign vec_sm_bitsReq_2_luma_inv[89] =87;
assign vec_sm_bitsReq_2_luma_inv[90] =140;
assign vec_sm_bitsReq_2_luma_inv[91] =200;
assign vec_sm_bitsReq_2_luma_inv[92] =117;
assign vec_sm_bitsReq_2_luma_inv[93] =213;
assign vec_sm_bitsReq_2_luma_inv[94] =176;
assign vec_sm_bitsReq_2_luma_inv[95] =224;
assign vec_sm_bitsReq_2_luma_inv[96] =131;
assign vec_sm_bitsReq_2_luma_inv[97] =44;
assign vec_sm_bitsReq_2_luma_inv[98] =194;
assign vec_sm_bitsReq_2_luma_inv[99] =56;
assign vec_sm_bitsReq_2_luma_inv[100] =39;
assign vec_sm_bitsReq_2_luma_inv[101] =138;
assign vec_sm_bitsReq_2_luma_inv[102] =27;
assign vec_sm_bitsReq_2_luma_inv[103] =42;
assign vec_sm_bitsReq_2_luma_inv[104] =201;
assign vec_sm_bitsReq_2_luma_inv[105] =162;
assign vec_sm_bitsReq_2_luma_inv[106] =78;
assign vec_sm_bitsReq_2_luma_inv[107] =168;
assign vec_sm_bitsReq_2_luma_inv[108] =141;
assign vec_sm_bitsReq_2_luma_inv[109] =30;
assign vec_sm_bitsReq_2_luma_inv[110] =75;
assign vec_sm_bitsReq_2_luma_inv[111] =106;
assign vec_sm_bitsReq_2_luma_inv[112] =114;
assign vec_sm_bitsReq_2_luma_inv[113] =54;
assign vec_sm_bitsReq_2_luma_inv[114] =156;
assign vec_sm_bitsReq_2_luma_inv[115] =99;
assign vec_sm_bitsReq_2_luma_inv[116] =166;
assign vec_sm_bitsReq_2_luma_inv[117] =154;
assign vec_sm_bitsReq_2_luma_inv[118] =216;
assign vec_sm_bitsReq_2_luma_inv[119] =169;
assign vec_sm_bitsReq_2_luma_inv[120] =15;
assign vec_sm_bitsReq_2_luma_inv[121] =198;
assign vec_sm_bitsReq_2_luma_inv[122] =177;
assign vec_sm_bitsReq_2_luma_inv[123] =170;
assign vec_sm_bitsReq_2_luma_inv[124] =210;
assign vec_sm_bitsReq_2_luma_inv[125] =45;
assign vec_sm_bitsReq_2_luma_inv[126] =57;
assign vec_sm_bitsReq_2_luma_inv[127] =217;
assign vec_sm_bitsReq_2_luma_inv[128] =108;
assign vec_sm_bitsReq_2_luma_inv[129] =228;
assign vec_sm_bitsReq_2_luma_inv[130] =204;
assign vec_sm_bitsReq_2_luma_inv[131] =103;
assign vec_sm_bitsReq_2_luma_inv[132] =147;
assign vec_sm_bitsReq_2_luma_inv[133] =120;
assign vec_sm_bitsReq_2_luma_inv[134] =135;
assign vec_sm_bitsReq_2_luma_inv[135] =51;
assign vec_sm_bitsReq_2_luma_inv[136] =91;
assign vec_sm_bitsReq_2_luma_inv[137] =225;
assign vec_sm_bitsReq_2_luma_inv[138] =180;
assign vec_sm_bitsReq_2_luma_inv[139] =94;
assign vec_sm_bitsReq_2_luma_inv[140] =157;
assign vec_sm_bitsReq_2_luma_inv[141] =151;
assign vec_sm_bitsReq_2_luma_inv[142] =229;
assign vec_sm_bitsReq_2_luma_inv[143] =121;
assign vec_sm_bitsReq_2_luma_inv[144] =118;
assign vec_sm_bitsReq_2_luma_inv[145] =109;
assign vec_sm_bitsReq_2_luma_inv[146] =181;
assign vec_sm_bitsReq_2_luma_inv[147] =240;
assign vec_sm_bitsReq_2_luma_inv[148] =214;
assign vec_sm_bitsReq_2_luma_inv[149] =195;
assign vec_sm_bitsReq_2_luma_inv[150] =79;
assign vec_sm_bitsReq_2_luma_inv[151] =60;
assign vec_sm_bitsReq_2_luma_inv[152] =205;
assign vec_sm_bitsReq_2_luma_inv[153] =55;
assign vec_sm_bitsReq_2_luma_inv[154] =31;
assign vec_sm_bitsReq_2_luma_inv[155] =220;
assign vec_sm_bitsReq_2_luma_inv[156] =43;
assign vec_sm_bitsReq_2_luma_inv[157] =115;
assign vec_sm_bitsReq_2_luma_inv[158] =119;
assign vec_sm_bitsReq_2_luma_inv[159] =142;
assign vec_sm_bitsReq_2_luma_inv[160] =163;
assign vec_sm_bitsReq_2_luma_inv[161] =178;
assign vec_sm_bitsReq_2_luma_inv[162] =221;
assign vec_sm_bitsReq_2_luma_inv[163] =139;
assign vec_sm_bitsReq_2_luma_inv[164] =202;
assign vec_sm_bitsReq_2_luma_inv[165] =107;
assign vec_sm_bitsReq_2_luma_inv[166] =232;
assign vec_sm_bitsReq_2_luma_inv[167] =58;
assign vec_sm_bitsReq_2_luma_inv[168] =244;
assign vec_sm_bitsReq_2_luma_inv[169] =199;
assign vec_sm_bitsReq_2_luma_inv[170] =158;
assign vec_sm_bitsReq_2_luma_inv[171] =46;
assign vec_sm_bitsReq_2_luma_inv[172] =155;
assign vec_sm_bitsReq_2_luma_inv[173] =241;
assign vec_sm_bitsReq_2_luma_inv[174] =95;
assign vec_sm_bitsReq_2_luma_inv[175] =184;
assign vec_sm_bitsReq_2_luma_inv[176] =172;
assign vec_sm_bitsReq_2_luma_inv[177] =226;
assign vec_sm_bitsReq_2_luma_inv[178] =122;
assign vec_sm_bitsReq_2_luma_inv[179] =124;
assign vec_sm_bitsReq_2_luma_inv[180] =61;
assign vec_sm_bitsReq_2_luma_inv[181] =211;
assign vec_sm_bitsReq_2_luma_inv[182] =182;
assign vec_sm_bitsReq_2_luma_inv[183] =233;
assign vec_sm_bitsReq_2_luma_inv[184] =245;
assign vec_sm_bitsReq_2_luma_inv[185] =185;
assign vec_sm_bitsReq_2_luma_inv[186] =173;
assign vec_sm_bitsReq_2_luma_inv[187] =110;
assign vec_sm_bitsReq_2_luma_inv[188] =167;
assign vec_sm_bitsReq_2_luma_inv[189] =218;
assign vec_sm_bitsReq_2_luma_inv[190] =230;
assign vec_sm_bitsReq_2_luma_inv[191] =215;
assign vec_sm_bitsReq_2_luma_inv[192] =125;
assign vec_sm_bitsReq_2_luma_inv[193] =47;
assign vec_sm_bitsReq_2_luma_inv[194] =186;
assign vec_sm_bitsReq_2_luma_inv[195] =174;
assign vec_sm_bitsReq_2_luma_inv[196] =206;
assign vec_sm_bitsReq_2_luma_inv[197] =143;
assign vec_sm_bitsReq_2_luma_inv[198] =171;
assign vec_sm_bitsReq_2_luma_inv[199] =203;
assign vec_sm_bitsReq_2_luma_inv[200] =234;
assign vec_sm_bitsReq_2_luma_inv[201] =111;
assign vec_sm_bitsReq_2_luma_inv[202] =179;
assign vec_sm_bitsReq_2_luma_inv[203] =59;
assign vec_sm_bitsReq_2_luma_inv[204] =62;
assign vec_sm_bitsReq_2_luma_inv[205] =246;
assign vec_sm_bitsReq_2_luma_inv[206] =236;
assign vec_sm_bitsReq_2_luma_inv[207] =242;
assign vec_sm_bitsReq_2_luma_inv[208] =222;
assign vec_sm_bitsReq_2_luma_inv[209] =237;
assign vec_sm_bitsReq_2_luma_inv[210] =183;
assign vec_sm_bitsReq_2_luma_inv[211] =126;
assign vec_sm_bitsReq_2_luma_inv[212] =248;
assign vec_sm_bitsReq_2_luma_inv[213] =123;
assign vec_sm_bitsReq_2_luma_inv[214] =249;
assign vec_sm_bitsReq_2_luma_inv[215] =231;
assign vec_sm_bitsReq_2_luma_inv[216] =159;
assign vec_sm_bitsReq_2_luma_inv[217] =219;
assign vec_sm_bitsReq_2_luma_inv[218] =227;
assign vec_sm_bitsReq_2_luma_inv[219] =188;
assign vec_sm_bitsReq_2_luma_inv[220] =189;
assign vec_sm_bitsReq_2_luma_inv[221] =187;
assign vec_sm_bitsReq_2_luma_inv[222] =250;
assign vec_sm_bitsReq_2_luma_inv[223] =63;
assign vec_sm_bitsReq_2_luma_inv[224] =207;
assign vec_sm_bitsReq_2_luma_inv[225] =175;
assign vec_sm_bitsReq_2_luma_inv[226] =223;
assign vec_sm_bitsReq_2_luma_inv[227] =238;
assign vec_sm_bitsReq_2_luma_inv[228] =247;
assign vec_sm_bitsReq_2_luma_inv[229] =235;
assign vec_sm_bitsReq_2_luma_inv[230] =253;
assign vec_sm_bitsReq_2_luma_inv[231] =127;
assign vec_sm_bitsReq_2_luma_inv[232] =252;
assign vec_sm_bitsReq_2_luma_inv[233] =190;
assign vec_sm_bitsReq_2_luma_inv[234] =243;
assign vec_sm_bitsReq_2_luma_inv[235] =239;
assign vec_sm_bitsReq_2_luma_inv[236] =191;
assign vec_sm_bitsReq_2_luma_inv[237] =254;
assign vec_sm_bitsReq_2_luma_inv[238] =255;
assign vec_sm_bitsReq_2_luma_inv[239] =251;
assign vec_sm_bitsReq_2_luma_inv[240] =85;
assign vec_sm_bitsReq_2_luma_inv[241] =21;
assign vec_sm_bitsReq_2_luma_inv[242] =69;
assign vec_sm_bitsReq_2_luma_inv[243] =5;
assign vec_sm_bitsReq_2_luma_inv[244] =81;
assign vec_sm_bitsReq_2_luma_inv[245] =17;
assign vec_sm_bitsReq_2_luma_inv[246] =65;
assign vec_sm_bitsReq_2_luma_inv[247] =1;
assign vec_sm_bitsReq_2_luma_inv[248] =84;
assign vec_sm_bitsReq_2_luma_inv[249] =20;
assign vec_sm_bitsReq_2_luma_inv[250] =68;
assign vec_sm_bitsReq_2_luma_inv[251] =4;
assign vec_sm_bitsReq_2_luma_inv[252] =80;
assign vec_sm_bitsReq_2_luma_inv[253] =16;
assign vec_sm_bitsReq_2_luma_inv[254] =64;
assign vec_sm_bitsReq_2_luma_inv[255] =0;

assign vec_sm_bitsReq_2_chroma_inv[0] =2;
assign vec_sm_bitsReq_2_chroma_inv[1] =8;
assign vec_sm_bitsReq_2_chroma_inv[2] =128;
assign vec_sm_bitsReq_2_chroma_inv[3] =32;
assign vec_sm_bitsReq_2_chroma_inv[4] =6;
assign vec_sm_bitsReq_2_chroma_inv[5] =9;
assign vec_sm_bitsReq_2_chroma_inv[6] =18;
assign vec_sm_bitsReq_2_chroma_inv[7] =72;
assign vec_sm_bitsReq_2_chroma_inv[8] =96;
assign vec_sm_bitsReq_2_chroma_inv[9] =144;
assign vec_sm_bitsReq_2_chroma_inv[10] =33;
assign vec_sm_bitsReq_2_chroma_inv[11] =132;
assign vec_sm_bitsReq_2_chroma_inv[12] =10;
assign vec_sm_bitsReq_2_chroma_inv[13] =24;
assign vec_sm_bitsReq_2_chroma_inv[14] =66;
assign vec_sm_bitsReq_2_chroma_inv[15] =129;
assign vec_sm_bitsReq_2_chroma_inv[16] =22;
assign vec_sm_bitsReq_2_chroma_inv[17] =36;
assign vec_sm_bitsReq_2_chroma_inv[18] =73;
assign vec_sm_bitsReq_2_chroma_inv[19] =160;
assign vec_sm_bitsReq_2_chroma_inv[20] =25;
assign vec_sm_bitsReq_2_chroma_inv[21] =70;
assign vec_sm_bitsReq_2_chroma_inv[22] =97;
assign vec_sm_bitsReq_2_chroma_inv[23] =82;
assign vec_sm_bitsReq_2_chroma_inv[24] =88;
assign vec_sm_bitsReq_2_chroma_inv[25] =148;
assign vec_sm_bitsReq_2_chroma_inv[26] =86;
assign vec_sm_bitsReq_2_chroma_inv[27] =37;
assign vec_sm_bitsReq_2_chroma_inv[28] =89;
assign vec_sm_bitsReq_2_chroma_inv[29] =12;
assign vec_sm_bitsReq_2_chroma_inv[30] =3;
assign vec_sm_bitsReq_2_chroma_inv[31] =133;
assign vec_sm_bitsReq_2_chroma_inv[32] =100;
assign vec_sm_bitsReq_2_chroma_inv[33] =145;
assign vec_sm_bitsReq_2_chroma_inv[34] =34;
assign vec_sm_bitsReq_2_chroma_inv[35] =101;
assign vec_sm_bitsReq_2_chroma_inv[36] =149;
assign vec_sm_bitsReq_2_chroma_inv[37] =136;
assign vec_sm_bitsReq_2_chroma_inv[38] =90;
assign vec_sm_bitsReq_2_chroma_inv[39] =192;
assign vec_sm_bitsReq_2_chroma_inv[40] =48;
assign vec_sm_bitsReq_2_chroma_inv[41] =165;
assign vec_sm_bitsReq_2_chroma_inv[42] =74;
assign vec_sm_bitsReq_2_chroma_inv[43] =7;
assign vec_sm_bitsReq_2_chroma_inv[44] =26;
assign vec_sm_bitsReq_2_chroma_inv[45] =13;
assign vec_sm_bitsReq_2_chroma_inv[46] =19;
assign vec_sm_bitsReq_2_chroma_inv[47] =76;
assign vec_sm_bitsReq_2_chroma_inv[48] =15;
assign vec_sm_bitsReq_2_chroma_inv[49] =112;
assign vec_sm_bitsReq_2_chroma_inv[50] =102;
assign vec_sm_bitsReq_2_chroma_inv[51] =153;
assign vec_sm_bitsReq_2_chroma_inv[52] =196;
assign vec_sm_bitsReq_2_chroma_inv[53] =161;
assign vec_sm_bitsReq_2_chroma_inv[54] =49;
assign vec_sm_bitsReq_2_chroma_inv[55] =98;
assign vec_sm_bitsReq_2_chroma_inv[56] =130;
assign vec_sm_bitsReq_2_chroma_inv[57] =164;
assign vec_sm_bitsReq_2_chroma_inv[58] =208;
assign vec_sm_bitsReq_2_chroma_inv[59] =38;
assign vec_sm_bitsReq_2_chroma_inv[60] =137;
assign vec_sm_bitsReq_2_chroma_inv[61] =40;
assign vec_sm_bitsReq_2_chroma_inv[62] =67;
assign vec_sm_bitsReq_2_chroma_inv[63] =28;
assign vec_sm_bitsReq_2_chroma_inv[64] =11;
assign vec_sm_bitsReq_2_chroma_inv[65] =152;
assign vec_sm_bitsReq_2_chroma_inv[66] =14;
assign vec_sm_bitsReq_2_chroma_inv[67] =23;
assign vec_sm_bitsReq_2_chroma_inv[68] =41;
assign vec_sm_bitsReq_2_chroma_inv[69] =134;
assign vec_sm_bitsReq_2_chroma_inv[70] =193;
assign vec_sm_bitsReq_2_chroma_inv[71] =77;
assign vec_sm_bitsReq_2_chroma_inv[72] =52;
assign vec_sm_bitsReq_2_chroma_inv[73] =240;
assign vec_sm_bitsReq_2_chroma_inv[74] =104;
assign vec_sm_bitsReq_2_chroma_inv[75] =224;
assign vec_sm_bitsReq_2_chroma_inv[76] =150;
assign vec_sm_bitsReq_2_chroma_inv[77] =71;
assign vec_sm_bitsReq_2_chroma_inv[78] =146;
assign vec_sm_bitsReq_2_chroma_inv[79] =29;
assign vec_sm_bitsReq_2_chroma_inv[80] =83;
assign vec_sm_bitsReq_2_chroma_inv[81] =170;
assign vec_sm_bitsReq_2_chroma_inv[82] =105;
assign vec_sm_bitsReq_2_chroma_inv[83] =92;
assign vec_sm_bitsReq_2_chroma_inv[84] =176;
assign vec_sm_bitsReq_2_chroma_inv[85] =35;
assign vec_sm_bitsReq_2_chroma_inv[86] =113;
assign vec_sm_bitsReq_2_chroma_inv[87] =87;
assign vec_sm_bitsReq_2_chroma_inv[88] =197;
assign vec_sm_bitsReq_2_chroma_inv[89] =53;
assign vec_sm_bitsReq_2_chroma_inv[90] =209;
assign vec_sm_bitsReq_2_chroma_inv[91] =212;
assign vec_sm_bitsReq_2_chroma_inv[92] =200;
assign vec_sm_bitsReq_2_chroma_inv[93] =93;
assign vec_sm_bitsReq_2_chroma_inv[94] =95;
assign vec_sm_bitsReq_2_chroma_inv[95] =50;
assign vec_sm_bitsReq_2_chroma_inv[96] =140;
assign vec_sm_bitsReq_2_chroma_inv[97] =116;
assign vec_sm_bitsReq_2_chroma_inv[98] =154;
assign vec_sm_bitsReq_2_chroma_inv[99] =106;
assign vec_sm_bitsReq_2_chroma_inv[100] =117;
assign vec_sm_bitsReq_2_chroma_inv[101] =166;
assign vec_sm_bitsReq_2_chroma_inv[102] =94;
assign vec_sm_bitsReq_2_chroma_inv[103] =169;
assign vec_sm_bitsReq_2_chroma_inv[104] =245;
assign vec_sm_bitsReq_2_chroma_inv[105] =213;
assign vec_sm_bitsReq_2_chroma_inv[106] =91;
assign vec_sm_bitsReq_2_chroma_inv[107] =51;
assign vec_sm_bitsReq_2_chroma_inv[108] =27;
assign vec_sm_bitsReq_2_chroma_inv[109] =30;
assign vec_sm_bitsReq_2_chroma_inv[110] =78;
assign vec_sm_bitsReq_2_chroma_inv[111] =138;
assign vec_sm_bitsReq_2_chroma_inv[112] =39;
assign vec_sm_bitsReq_2_chroma_inv[113] =75;
assign vec_sm_bitsReq_2_chroma_inv[114] =42;
assign vec_sm_bitsReq_2_chroma_inv[115] =204;
assign vec_sm_bitsReq_2_chroma_inv[116] =229;
assign vec_sm_bitsReq_2_chroma_inv[117] =141;
assign vec_sm_bitsReq_2_chroma_inv[118] =168;
assign vec_sm_bitsReq_2_chroma_inv[119] =99;
assign vec_sm_bitsReq_2_chroma_inv[120] =162;
assign vec_sm_bitsReq_2_chroma_inv[121] =114;
assign vec_sm_bitsReq_2_chroma_inv[122] =103;
assign vec_sm_bitsReq_2_chroma_inv[123] =177;
assign vec_sm_bitsReq_2_chroma_inv[124] =31;
assign vec_sm_bitsReq_2_chroma_inv[125] =225;
assign vec_sm_bitsReq_2_chroma_inv[126] =54;
assign vec_sm_bitsReq_2_chroma_inv[127] =181;
assign vec_sm_bitsReq_2_chroma_inv[128] =157;
assign vec_sm_bitsReq_2_chroma_inv[129] =201;
assign vec_sm_bitsReq_2_chroma_inv[130] =228;
assign vec_sm_bitsReq_2_chroma_inv[131] =216;
assign vec_sm_bitsReq_2_chroma_inv[132] =156;
assign vec_sm_bitsReq_2_chroma_inv[133] =118;
assign vec_sm_bitsReq_2_chroma_inv[134] =79;
assign vec_sm_bitsReq_2_chroma_inv[135] =180;
assign vec_sm_bitsReq_2_chroma_inv[136] =194;
assign vec_sm_bitsReq_2_chroma_inv[137] =56;
assign vec_sm_bitsReq_2_chroma_inv[138] =131;
assign vec_sm_bitsReq_2_chroma_inv[139] =217;
assign vec_sm_bitsReq_2_chroma_inv[140] =44;
assign vec_sm_bitsReq_2_chroma_inv[141] =244;
assign vec_sm_bitsReq_2_chroma_inv[142] =158;
assign vec_sm_bitsReq_2_chroma_inv[143] =210;
assign vec_sm_bitsReq_2_chroma_inv[144] =57;
assign vec_sm_bitsReq_2_chroma_inv[145] =108;
assign vec_sm_bitsReq_2_chroma_inv[146] =45;
assign vec_sm_bitsReq_2_chroma_inv[147] =175;
assign vec_sm_bitsReq_2_chroma_inv[148] =147;
assign vec_sm_bitsReq_2_chroma_inv[149] =109;
assign vec_sm_bitsReq_2_chroma_inv[150] =241;
assign vec_sm_bitsReq_2_chroma_inv[151] =135;
assign vec_sm_bitsReq_2_chroma_inv[152] =198;
assign vec_sm_bitsReq_2_chroma_inv[153] =151;
assign vec_sm_bitsReq_2_chroma_inv[154] =119;
assign vec_sm_bitsReq_2_chroma_inv[155] =120;
assign vec_sm_bitsReq_2_chroma_inv[156] =214;
assign vec_sm_bitsReq_2_chroma_inv[157] =107;
assign vec_sm_bitsReq_2_chroma_inv[158] =121;
assign vec_sm_bitsReq_2_chroma_inv[159] =250;
assign vec_sm_bitsReq_2_chroma_inv[160] =233;
assign vec_sm_bitsReq_2_chroma_inv[161] =142;
assign vec_sm_bitsReq_2_chroma_inv[162] =182;
assign vec_sm_bitsReq_2_chroma_inv[163] =221;
assign vec_sm_bitsReq_2_chroma_inv[164] =55;
assign vec_sm_bitsReq_2_chroma_inv[165] =220;
assign vec_sm_bitsReq_2_chroma_inv[166] =43;
assign vec_sm_bitsReq_2_chroma_inv[167] =255;
assign vec_sm_bitsReq_2_chroma_inv[168] =115;
assign vec_sm_bitsReq_2_chroma_inv[169] =171;
assign vec_sm_bitsReq_2_chroma_inv[170] =155;
assign vec_sm_bitsReq_2_chroma_inv[171] =110;
assign vec_sm_bitsReq_2_chroma_inv[172] =205;
assign vec_sm_bitsReq_2_chroma_inv[173] =186;
assign vec_sm_bitsReq_2_chroma_inv[174] =173;
assign vec_sm_bitsReq_2_chroma_inv[175] =122;
assign vec_sm_bitsReq_2_chroma_inv[176] =202;
assign vec_sm_bitsReq_2_chroma_inv[177] =218;
assign vec_sm_bitsReq_2_chroma_inv[178] =58;
assign vec_sm_bitsReq_2_chroma_inv[179] =230;
assign vec_sm_bitsReq_2_chroma_inv[180] =46;
assign vec_sm_bitsReq_2_chroma_inv[181] =174;
assign vec_sm_bitsReq_2_chroma_inv[182] =195;
assign vec_sm_bitsReq_2_chroma_inv[183] =167;
assign vec_sm_bitsReq_2_chroma_inv[184] =139;
assign vec_sm_bitsReq_2_chroma_inv[185] =178;
assign vec_sm_bitsReq_2_chroma_inv[186] =185;
assign vec_sm_bitsReq_2_chroma_inv[187] =232;
assign vec_sm_bitsReq_2_chroma_inv[188] =111;
assign vec_sm_bitsReq_2_chroma_inv[189] =60;
assign vec_sm_bitsReq_2_chroma_inv[190] =234;
assign vec_sm_bitsReq_2_chroma_inv[191] =159;
assign vec_sm_bitsReq_2_chroma_inv[192] =226;
assign vec_sm_bitsReq_2_chroma_inv[193] =246;
assign vec_sm_bitsReq_2_chroma_inv[194] =184;
assign vec_sm_bitsReq_2_chroma_inv[195] =211;
assign vec_sm_bitsReq_2_chroma_inv[196] =163;
assign vec_sm_bitsReq_2_chroma_inv[197] =61;
assign vec_sm_bitsReq_2_chroma_inv[198] =123;
assign vec_sm_bitsReq_2_chroma_inv[199] =172;
assign vec_sm_bitsReq_2_chroma_inv[200] =187;
assign vec_sm_bitsReq_2_chroma_inv[201] =238;
assign vec_sm_bitsReq_2_chroma_inv[202] =249;
assign vec_sm_bitsReq_2_chroma_inv[203] =125;
assign vec_sm_bitsReq_2_chroma_inv[204] =183;
assign vec_sm_bitsReq_2_chroma_inv[205] =47;
assign vec_sm_bitsReq_2_chroma_inv[206] =143;
assign vec_sm_bitsReq_2_chroma_inv[207] =199;
assign vec_sm_bitsReq_2_chroma_inv[208] =179;
assign vec_sm_bitsReq_2_chroma_inv[209] =248;
assign vec_sm_bitsReq_2_chroma_inv[210] =124;
assign vec_sm_bitsReq_2_chroma_inv[211] =206;
assign vec_sm_bitsReq_2_chroma_inv[212] =237;
assign vec_sm_bitsReq_2_chroma_inv[213] =59;
assign vec_sm_bitsReq_2_chroma_inv[214] =239;
assign vec_sm_bitsReq_2_chroma_inv[215] =126;
assign vec_sm_bitsReq_2_chroma_inv[216] =215;
assign vec_sm_bitsReq_2_chroma_inv[217] =222;
assign vec_sm_bitsReq_2_chroma_inv[218] =251;
assign vec_sm_bitsReq_2_chroma_inv[219] =189;
assign vec_sm_bitsReq_2_chroma_inv[220] =62;
assign vec_sm_bitsReq_2_chroma_inv[221] =219;
assign vec_sm_bitsReq_2_chroma_inv[222] =254;
assign vec_sm_bitsReq_2_chroma_inv[223] =191;
assign vec_sm_bitsReq_2_chroma_inv[224] =203;
assign vec_sm_bitsReq_2_chroma_inv[225] =242;
assign vec_sm_bitsReq_2_chroma_inv[226] =231;
assign vec_sm_bitsReq_2_chroma_inv[227] =190;
assign vec_sm_bitsReq_2_chroma_inv[228] =127;
assign vec_sm_bitsReq_2_chroma_inv[229] =235;
assign vec_sm_bitsReq_2_chroma_inv[230] =236;
assign vec_sm_bitsReq_2_chroma_inv[231] =188;
assign vec_sm_bitsReq_2_chroma_inv[232] =253;
assign vec_sm_bitsReq_2_chroma_inv[233] =243;
assign vec_sm_bitsReq_2_chroma_inv[234] =227;
assign vec_sm_bitsReq_2_chroma_inv[235] =207;
assign vec_sm_bitsReq_2_chroma_inv[236] =63;
assign vec_sm_bitsReq_2_chroma_inv[237] =247;
assign vec_sm_bitsReq_2_chroma_inv[238] =223;
assign vec_sm_bitsReq_2_chroma_inv[239] =252;
assign vec_sm_bitsReq_2_chroma_inv[240] =85;
assign vec_sm_bitsReq_2_chroma_inv[241] =21;
assign vec_sm_bitsReq_2_chroma_inv[242] =69;
assign vec_sm_bitsReq_2_chroma_inv[243] =5;
assign vec_sm_bitsReq_2_chroma_inv[244] =81;
assign vec_sm_bitsReq_2_chroma_inv[245] =17;
assign vec_sm_bitsReq_2_chroma_inv[246] =65;
assign vec_sm_bitsReq_2_chroma_inv[247] =1;
assign vec_sm_bitsReq_2_chroma_inv[248] =84;
assign vec_sm_bitsReq_2_chroma_inv[249] =20;
assign vec_sm_bitsReq_2_chroma_inv[250] =68;
assign vec_sm_bitsReq_2_chroma_inv[251] =4;
assign vec_sm_bitsReq_2_chroma_inv[252] =80;
assign vec_sm_bitsReq_2_chroma_inv[253] =16;
assign vec_sm_bitsReq_2_chroma_inv[254] =64;
assign vec_sm_bitsReq_2_chroma_inv[255] =0;

endmodule


