module decBpvBlock #(parameter ssm_idx = 0)
(

  input mode_BP,
  input use2x2,
  input [127:0] suffix,
  output [7:0]  bpv_size
);



endmodule
